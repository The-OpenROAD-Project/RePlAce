../library/nangate45/NangateOpenCellLibrary.lef